module mux4to1_str_tb;
reg [0:3]I;
reg [1:0]S;
wire Y;

mux4to1_str dut(.I(I), .S(S), .Y(Y));

initial
begin
    I = 4'b1010;
    S = 2'b00;
    #100
    I = 4'b1010;
    S = 2'b01;
    #100
    I = 4'b1010;
    S = 2'b10;
    #100 
    I = 4'b1010;
    S = 2'b11;
 end
 endmodule
